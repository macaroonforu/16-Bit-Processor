module proc(DIN, Resetn, Clock, Run, DOUT, ADDR, W);
    parameter N = 3; 
	input [15:0] DIN;
    input Resetn, Clock, Run;
    output wire [15:0] DOUT;
    output wire [15:0] ADDR;
    output wire W;

    wire [0:7] R_in; // r0, ..., r7 register enables
    reg rX_in, IR_in, ADDR_in, Done, DOUT_in, A_in, G_in, AddSub, ALU_and, F_in;
    reg [2:0] Tstep_Q, Tstep_D;
    reg [15:0] BusWires;
    reg [3:0] Select; // BusWires selector
    reg [16:0] Sum;
    wire [2:0] III, rX, rY; // instruction opcode and register operands
    wire [15:0] r0, r1, r2, r3, r4, r5, r6, pc, A;
    wire [15:0] G;
    wire [15:0] IR;
    reg pc_incr;    // used to increment the pc
    reg pc_in;      // used to load the pc
	reg lr_in; //used to load the lr
    reg W_D;        // used for write signal
	reg do_shift; 
    wire Imm;
	reg sp_incr; 
	reg sp_decr; 
	wire [15:0] sp; 
   
   
    assign III = IR[15:13];
    assign rX = IR[11:9];
    assign rY = IR[2:0];
	assign Imm = IR[12];
	
	
	wire d; 
	assign d = IR[7]; 
	
	wire[5:0] cmpShift; 
	assign cmpShift = IR[8:3];
	
	wire[1:0] shift_type; 
	assign shift_type = IR[6:5];
	
    dec3to8 decX (rX_in, rX, R_in); // produce r0 - r7 register enables
	
	wire [2:0] concat; 
    parameter T0 = 3'b000, T1 = 3'b001, T2 = 3'b010, T3 = 3'b011, T4 = 3'b100, T5 = 3'b101;
    // Control FSM state table
    always @(Tstep_Q, Run, Done)
        case (Tstep_Q)
            T0: // instruction fetch
                if (~Run) Tstep_D = T0;
                else Tstep_D = T1;
            T1: // wait cycle for synchronous memory
                Tstep_D = T2;
            T2: // this time step stores the instruction word in IR
                Tstep_D = T3;
            T3: if (Done) Tstep_D = T0;
                else Tstep_D = T4;
            T4: if (Done) Tstep_D = T0;
                else Tstep_D = T5;
            T5: // instructions end after this time step
                Tstep_D = T0;
            default: Tstep_D = 3'bxxx;
        endcase

    /* OPCODE format: III M XXX DDDDDDDDD, where 
    *     III = instruction, M = Immediate, XXX = rX. If M = 0, DDDDDDDDD = 000000YYY = rY
    *     If M = 1, DDDDDDDDD = #D is the immediate operand 
    *
    *  III M  Instruction   Description
    *  --- -  -----------   -----------
    *  000 0: mv   rX,rY    rX <- rY
    *  000 1: mv   rX,#D    rX <- D (sign extended)
    *  001 1: mvt  rX,#D    rX <- D << 8
    *  010 0: add  rX,rY    rX <- rX + rY
    *  010 1: add  rX,#D    rX <- rX + D
    *  011 0: sub  rX,rY    rX <- rX - rY
    *  011 1: sub  rX,#D    rX <- rX - D
    *  100 0: ld   rX,[rY]  rX <- [rY]
    *  101 0: st   rX,[rY]  [rY] <- rX
	
	
    *  110 0: and  rX,rY    rX <- rX & rY
    *  110 1: and  rX,#D    rX <- rX & D 
	
	
	*  100 1: pop  rX       rX <- [sp], sp<- sp+1 
	   101 1: push rX       sp<- sp-1, [sp] <- rX 
	   
	   
	   111 0: cmp  rX, rY   performs rX-rY, sets flags
	   111 1: cmp  rX, #D   performs rX - D, sets flags 
			  */
	
    parameter mv = 3'b000, mvt = 3'b001, add = 3'b010, sub = 3'b011, ld = 3'b100, st = 3'b101,
	     and_ = 3'b110, pop = 3'b100, push = 3'b101, cmp = 3'b111; 
		 
    // selectors for the BusWires multiplexer
    parameter _R0 = 4'b0000, _R1 = 4'b0001, _R2 = 4'b0010, _R3 = 4'b0011, _R4 = 4'b0100,
        _R5 = 4'b0101, _R6 = 4'b0110, _PC = 4'b0111, _G = 4'b1000, 
        _IR8_IR8_0 /* signed-extended immediate data */ = 4'b1001, 
        _IR7_0_0 /* immediate data << 8 */ = 4'b1010,
        _DIN /* data-in from memory */ = 4'b1011, 
		_SHIFT_IR8 = 4'b1100; 
		
    // Control FSM outputs
    always @(*) begin
        // default values for control signals
        rX_in = 1'b0; A_in = 1'b0; G_in = 1'b0; IR_in = 1'b0; DOUT_in = 1'b0; ADDR_in = 1'b0; 
        //Select = 4'bxxxx; 
		AddSub = 1'b0; ALU_and = 1'b0; W_D = 1'b0; Done = 1'b0;
        pc_in = R_in[7]; 
		lr_in = R_in[6]; 
		F_in = 1'b0; 

		/* default pc enable */pc_incr = 1'b0; sp_incr = 1'b0; sp_decr = 1'b0; do_shift = 1'b0;
		
        case (Tstep_Q)
            T0: begin // fetch the instruction
                Select = _PC;  //put pc onto the bus wires (same cycle) 
                ADDR_in = 1'b1; //Enable reg_adr to receive what is on the bus wires on the next clock cycle 
                pc_incr = Run; //pc_incr is the enable signal on the pc register that tells it to increment itself 
            end
            T1: begin //wait cycle for synchronous memory 
				//address now = pc 
				//WREN = 0, so it means that we will read from the address stored at the ADDR port
				//q <= data stored at pc 
				Select = _DIN; 
                //;
			end 
            T2: begin // store instruction on DIN in IR 
				//q is connected to DIN so when ir = 1, we are getting DIN
				//and DIN is what we read from pc's address in the memory unit 
				Select = _DIN; 
                IR_in = 1'b1; 
			end 
            T3: // define signals in T3
                case (III)
                    mv: begin
                        if (!Imm) Select = rY;            // mv rX, rY
                        else Select = _IR8_IR8_0;        // mv rX, #D
                        rX_in = 1'b1;                   // enable the rX register
                        Done = 1'b1;
                    end
                    mvt: begin
					
						if(Imm)begin //code for a move top 
                        Select = _IR7_0_0; 
						rX_in = 1'b1; 
						Done = 1'b1; 
						end 
						//concat[2]=c concat[1] = n concat[0] = z 
						else begin      //code for a b{cond}
						Select = _PC;  //Put the PC on the buswires 
						A_in = 1'b1;  //Put the PC in the A register 
						case(rX)     //IR[11:9] specifies the condition 
							/*B*/3'b000:  	Done = 0;     					 //always take the branch 
							/*BEQ*/3'b001:  Done = (concat[0]==1'b1)? 0:1;   //if z flag = 1, we have a zero condition, so continue on 
							/*BNE*/3'b010:  Done = (concat[0]==1'b0)? 0:1;  //If z flag = 0, we have a nonzero condition, so continue on 
							/*BCC*/3'b011:  Done = (concat[2]==1'b0)? 0:1;  //if c flag = 0, we have a carry clear condition 
							/*BCS*/3'b100:  Done = (concat[2]==1'b1)? 0:1; //if c flag = 1, we have a carry set condition 
							/*BPL*/3'b101:  Done = (concat[1]==1'b0)? 0:1; //if n flag = 0, we have a plus condition 
							/*BMI*/3'b110:  Done = (concat[1]==1'b1)? 0:1; //if n flag = 1, we have a minus condition  
							/*BL*/ 3'b111:  lr_in = 1'b1;  //load the lr (R6) with the pc's current value 
						endcase 
						end 
                    end
                    add, sub, and_: begin
                        Select = rX; 
						A_in = 1'b1; 	
                    end
                    ld: begin
						Select = rY;  //Put rY onto the Bus Wires 
						ADDR_in = 1'b1; //Enable the address register to receive what is on the bus wires in the next clock cycle 
						if(rY==3'b101)begin 
							sp_incr = 1'b1; //pop
						end 	
                    end
					
					st: begin 
						if(rY==3'b101)begin  
							sp_decr = 1'b1;  //push
						end 
						else begin 
							Select = rY;  //Put rY onto the Bus Wires 
							ADDR_in = 1'b1; //Enable the address register to receive what is on the bus wires in the next clock cycle 
						end 
						
					end 
					
					cmp: begin 
						Select = rX; 
						A_in = 1'b1;  //Take in rX 
					end 
					
                    default: ;
                endcase
            T4: // define signals T2
                case (III)
                    add: begin
                        Select = Imm? _IR8_IR8_0: rY;
						G_in = 1'b1; 
						F_in = 1'b1; 
						AddSub = 1'b0; 
                    end
                    sub: begin
                        Select = Imm? _IR8_IR8_0: rY;
						G_in = 1'b1; 
						F_in = 1'b1;
						AddSub = 1'b1; 
                    end
                    and_: begin
                        Select = Imm? _IR8_IR8_0: rY;
						G_in = 1'b1; 
						F_in = 1'b1;
						ALU_and = 1'b1; 
                    end
					mvt: begin   
						Select = _IR8_IR8_0; //Put the branch offset onto the bus Wires
						G_in = 1;  //ALU adds PC + branch offset in the same cycle and outputs that to G register 
						AddSub = 1'b0; 
					end 
                    ld: begin //Read the value from the address (rY) and output it to DIN 
						W_D = 1'b0; 
						
					end 
                    st: begin
					
						if(rY == 3'b101)begin 
							Select = rY;  //code for the push 
							ADDR_in = 1'b1; 
						end 
						
						else begin 
							Select = rX; //Put rX onto the bus Wires 
							DOUT_in = 1'b1; //Enable the data register to receive data from the bus wires on the next clock cycle (this data is rX) 
							W_D = 1'b1; //Write the value at Data port to the address at address port of memory (write data rx to address rY) 
							Done = 1'b1; 
						end 
                    end
					
					
					cmp: begin  
						if(Imm) begin  //cmp Rx, #D
							Select = _IR8_IR8_0; 
							AddSub = 1'b1; 
							F_in = 1'b1; 
							Done = 1'b1; 
						end 
						
						else begin 
							if(cmpShift == 6'b0)begin //cmp Rx, Ry 
								Select = rY; 
								AddSub = 1'b1; 
								F_in = 1'b1; 
								Done = 1'b1;
							end 
							
							else begin //Shift Rx, #D
								Select = d? _SHIFT_IR8: rY;// shift by amount DDDD or rY
								do_shift = 1'b1;
								G_in = 1'b1; 
								F_in = 1'b1;
							end
						end 
					end 
					
                    default: ; 
                endcase
            T5: // define T3
                case (III)
                    add, sub, and_: begin
                        Select = _G; 
						rX_in = 1'b1;
						Done = 1'b1; 
                    end
					
                    ld: begin
							Select = _DIN;  //Put DIN onto the bus Wires
							rX_in = 1'b1;  //Enable rX to recieve data on the bus Wires (the sum)in the following clock cycles 
							Done = 1'b1;  
                    end 
					
					st: begin 
						if(rY ==3'b101) begin //push 
							Select = rX;  //Put DIN onto the bus Wires
							DOUT_in = 1'b1;  //Enable rX to recieve data on the bus Wires (the sum)in the following clock cycles 
							Done = 1'b1;
							W_D = 1'b1; 
						end  
					end 
					
					mvt: begin 
						Select = _G;    //Put G on the BusWires (pc + branch offset) 
						pc_in = 1'b1;  //Pc takes in G so we now go to a new branch 
						Done = 1'b1; 
					end
					
					cmp: begin 
						Select = _G; 
						rX_in = 1'b1; 
						Done = 1'b1; 
					end 
					
                    default: ;
                endcase
            default: ;
        endcase
    end   
   
    // Control FSM flip-flops
    always @(posedge Clock)
        if (!Resetn)
            Tstep_Q <= T0;
        else
            Tstep_Q <= Tstep_D;   
   
    regn reg_0 (BusWires, Resetn, R_in[0], Clock, r0);
    regn reg_1 (BusWires, Resetn, R_in[1], Clock, r1);
    regn reg_2 (BusWires, Resetn, R_in[2], Clock, r2);
    regn reg_3 (BusWires, Resetn, R_in[3], Clock, r3);
    regn reg_4 (BusWires, Resetn, R_in[4], Clock, r4);
    // regn reg_5 (BusWires, Resetn, R_in[5], Clock, r5);
    regn lr (BusWires, Resetn, lr_in, Clock, r6);

    // r7 is program counter
    // module pc_count(R, Resetn, Clock, E, L, Q);
    pc_count reg_pc (BusWires, Resetn, Clock, pc_incr, pc_in, pc);
	
	sp_count reg_sp (BusWires, Resetn, Clock, sp_incr, sp_decr, R_in[5], r5); 

    regn reg_A (BusWires, Resetn, A_in, Clock, A);
    regn reg_DOUT (BusWires, Resetn, DOUT_in, Clock, DOUT);
    regn reg_ADDR (BusWires, Resetn, ADDR_in, Clock, ADDR);
    regn reg_IR (DIN, Resetn, IR_in, Clock, IR);
    flipflop reg_W (W_D, Resetn, Clock, W);
	
	//Condition Code stuff 
	regn #(.n(N)) cond_code({Sum[16], Sum[15], (Sum==17'b0)}, Resetn, F_in, Clock, concat); 
	
    // alu
    always @(*)
		if (!AddSub && !do_shift && !ALU_and)begin 
			Sum = A + BusWires; 
		end 
		
        else if (AddSub) begin 
			Sum = A + ~BusWires + 16'b1; 
		end
		
		else if (do_shift) begin  //A is Rx, BusWires is Op2 
			case (shift_type)
				2'b00: Sum = A << BusWires[3:0];  //LSL
				2'b01: Sum = A >> BusWires[3:0]; //LSR
				2'b10: Sum = {{16{A[15]}}, A} >> BusWires[3:0]; //ASR
				2'b11: Sum = (A>>BusWires[3:0])|(A<<(16'd16-BusWires[3:0])); //ROR
			endcase
		end
		
		else if (ALU_and) begin
			Sum = A & BusWires;
		end
		
    regn reg_G (Sum[15:0], Resetn, G_in, Clock, G);
	
    // define the internal processor bus
    always @(*)
        case (Select)
            _R0: BusWires = r0;
            _R1: BusWires = r1;
            _R2: BusWires = r2;
            _R3: BusWires = r3;
            _R4: BusWires = r4;
            _R5: BusWires = r5;
            _R6: BusWires = r6;
            _PC: BusWires = pc;
            _G: BusWires = G;
            _IR8_IR8_0: BusWires = {{7{IR[8]}}, IR[8:0]}; // sign extended
            _IR7_0_0: BusWires = {IR[7:0], 8'b0};
            _DIN: BusWires = DIN;
			_SHIFT_IR8: BusWires = {{12{IR[3]}}, IR[3:0]}; 
            default: BusWires = 16'bx;
        endcase
endmodule

module pc_count(R, Resetn, Clock, E, L, Q);
    input [15:0] R;
    input Resetn, Clock, E, L;
    output [15:0] Q;
    reg [15:0] Q;
   
    always @(posedge Clock)
        if (!Resetn)
            Q <= 16'b0;
        else if (L)
            Q <= R;
        else if (E)
            Q <= Q + 1'b1;
endmodule

module sp_count(R, Resetn, Clock, U, D, L, Q); 
	input [15:0] R; 
	input Resetn, Clock, U, D, L; 
	output [15:0] Q; 
	reg [15:0] Q; 
	
	always@(posedge Clock) 
		if(!Resetn)
			Q <= 16'b0; 
		else if (L) 
			Q <= R; 
		else if (U)
			Q <= Q + 1'b1; 
		else if (D) 
			Q <= Q - 1'b1;
endmodule 

module dec3to8(E, W, Y);
    input E; // enable
    input [2:0] W;
    output [0:7] Y;
    reg [0:7] Y;
   
    always @(*)
        if (E == 0)
            Y = 8'b00000000;
        else
            case (W)
                3'b000: Y = 8'b10000000;
                3'b001: Y = 8'b01000000;
                3'b010: Y = 8'b00100000;
                3'b011: Y = 8'b00010000;
                3'b100: Y = 8'b00001000;
                3'b101: Y = 8'b00000100;
                3'b110: Y = 8'b00000010;
                3'b111: Y = 8'b00000001;
            endcase
endmodule

module regn(R, Resetn, E, Clock, Q);
    parameter n = 16;
    input [n-1:0] R;
    input Resetn, E, Clock;
    output [n-1:0] Q;
    reg [n-1:0] Q;

    always @(posedge Clock)
        if (!Resetn)
            Q <= 0;
        else if (E)
            Q <= R;
endmodule
